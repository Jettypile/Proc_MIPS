/*
    CS/ECE 552 Spring '20
    Homework #1, Problem 2
    
    a 4-bit CLA module
*/
module cla_4b(A, B, C_in, S, C_out);

    // declare constant for size of inputs, outputs (N)
    parameter   N = 4;

    input [N-1: 0] A, B;
    input          C_in;
    output [N-1:0] S;
    output         C_out;

    // YOUR CODE HERE
    wire [3:0] g, p;
    genPropLogic gpblock0(.A(A), .B(B), .g(g), .p(p), .superG(), .superP());

    wire [3:0] sub_carry;
    claLogicBlock carryLogic(.G(g), .P(p), .C_in(C_in), .C_out(sub_carry));
    assign C_out = sub_carry[3];

    // SUM Calculation
    fullAdder_1b fa_sum0(.A(A[0]), .B(B[0]), .C_in(C_in), .S(S[0]), .C_out());
    fullAdder_1b fa_sum1(.A(A[1]), .B(B[1]), .C_in(sub_carry[0]), .S(S[1]), .C_out());
    fullAdder_1b fa_sum2(.A(A[2]), .B(B[2]), .C_in(sub_carry[1]), .S(S[2]), .C_out());
    fullAdder_1b fa_sum3(.A(A[3]), .B(B[3]), .C_in(sub_carry[2]), .S(S[3]), .C_out());

endmodule
